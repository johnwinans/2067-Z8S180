//**************************************************************************
//
//    Copyright (C) 2025  John Winans
//
//    This library is free software; you can redistribute it and/or
//    modify it under the terms of the GNU Lesser General Public
//    License as published by the Free Software Foundation; either
//    version 2.1 of the License, or (at your option) any later version.
//
//    This library is distributed in the hope that it will be useful,
//    but WITHOUT ANY WARRANTY; without even the implied warranty of
//    MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the GNU
//    Lesser General Public License for more details.
//
//    You should have received a copy of the GNU Lesser General Public
//    License along with this library; if not, write to the Free Software
//    Foundation, Inc., 51 Franklin Street, Fifth Floor, Boston, MA  02110-1301
//    USA
//
//**************************************************************************

`timescale 1ns/1ns
`default_nettype none

module tb ();

    reg     reset   = 0;
    reg     clk     = 0;
    wire    ay_clk;
    wire    noise_out;

    localparam CLK_FREQ         = 25000000;
    localparam CLK_PERIOD       = (1.0/CLK_FREQ)*1000000000;
    localparam AY_CLK_FREQ      = 1789773;
    localparam AY_CLK_PERIOD    = (1.0/AY_CLK_FREQ)*1000000000;

    wire [4:0] NOISE_PERIOD     = 9;

    always #(CLK_PERIOD/2) clk = ~clk;

    prescaler #(
        .IN_FREQ(CLK_FREQ),
        .OUT_FREQ(AY_CLK_FREQ)
    ) the_prescaler (
        .reset(reset),
        .clk(clk),
        .out(ay_clk)
    );

    ay_noise noise (
        .reset(reset),
        .clk(clk),
        .ay_clk(ay_clk),
        .period(NOISE_PERIOD),
        .out(noise_out)
    );

    initial begin
        $dumpfile( { `__FILE__, "cd" } );
        $dumpvars;

        #(CLK_PERIOD*4);
        reset <= 1;
        #(CLK_PERIOD*4);
        reset <= 0;
        #(CLK_PERIOD*4);

        //#(NOISE_PERIOD*AY_CLK_PERIOD*1000);
        #1000000;

        $finish;
    end

endmodule
